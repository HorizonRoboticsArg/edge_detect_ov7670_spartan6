--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package paquete_multiplexor is

type vector16x16bits is array (15 downto 0) of std_logic_vector(15 downto 0);

end paquete_multiplexor;

